../ips/axi/axi_demux.sv