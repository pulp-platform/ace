package ace_test_pkg;
`define _ACE_TEST_PKG
`include "ace/ace_beat_types.svh"
`include "ace/ace_driver.svh"
`include "ace/ace_monitor.svh"
`include "ace/ace_sequencer.svh"
`include "ace/ace_agent.svh"
endpackage