../ips/axi/axi_demux_simple.sv