package ccu_ctrl_pkg;

    typedef enum logic { MEMORY_UNIT, SNOOP_UNIT } dest_t;

endpackage