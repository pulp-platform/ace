package cache_test_pkg;
`define _CACHE_TEST_PKG
`include "cache/cache_top_agent.svh"
endpackage