../ips/axi/axi_mux.sv