package cache_test_pkg;
`define _CACHE_TEST_PKG
`include "cache/cache_beat_types.svh"
`include "cache/cache_sequencer.svh"
`include "cache/cache_scoreboard.svh"
`include "cache/cache_top_agent.svh"
endpackage