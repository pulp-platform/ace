../ips/axi/axi_cut.sv